module blowfish

struct CryptTest {
	key 	[]byte
	ins  	[]byte
	out 	[]byte
}

fn test_main() {
	rs := [
		CryptTest{
			key: [byte(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00]
			ins: [byte(0x00), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00]
			out: [byte(0x4E), 0xF9, 0x97, 0x45, 0x61, 0x98, 0xDD, 0x78]
		},
		CryptTest{
			key: [byte(0xFF), 0xFF, 0xFF, 0xFF, 0xFF, 0xFF, 0xFF, 0xFF]
			ins: [byte(0xFF), 0xFF, 0xFF, 0xFF, 0xFF, 0xFF, 0xFF, 0xFF]
			out: [byte(0x51), 0x86, 0x6F, 0xD5, 0xB8, 0x5E, 0xCB, 0x8A]
		},
		CryptTest{
			key: [byte(0x30), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x00]
			ins: [byte(0x10), 0x00, 0x00, 0x00, 0x00, 0x00, 0x00, 0x01]
			out: [byte(0x7D), 0x85, 0x6F, 0x9A, 0x61, 0x30, 0x63, 0xF2]
		}
	]

	for s in rs {
		c := blowfish.new_cipher(s.key) or {
			panic(err)
		}

		mut ct := []byte{len: s.out.len}
		c.encrypt(mut ct, s.ins)

		for j, v in ct {
			assert v == s.out[j]
		}
	}
}