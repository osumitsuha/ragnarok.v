module constants

pub enum Packets {
	osu_change_action = 0
    osu_send_public_message = 1
    osu_logout = 2
    osu_request_status_update = 3
    osu_ping = 4
    cho_user_id = 5
    cho_cmd_err = 6  
    cho_send_message = 7
    cho_pong = 8
    cho_handle_irc_change_username = 9
    cho_handle_irc_quit = 10  
    cho_user_stats = 11
    cho_user_logout = 12
    cho_spectator_joined = 13
    cho_spectator_left = 14
    cho_spectate_frames = 15
    osu_start_spectating = 16
    osu_stop_spectating = 17
    osu_spectate_frames = 18
    cho_version_update = 19
    osu_error_report = 20  
    osu_cant_spectate = 21
    cho_spectator_cant_spectate = 22
    cho_get_attention = 23
    cho_notification = 24
    osu_send_private_message = 25
    cho_update_match = 26
    cho_new_match = 27
    cho_dispose_match = 28
    osu_part_lobby = 29
    osu_join_lobby = 30
    osu_create_match = 31
    osu_join_match = 32
    osu_part_match = 33
    cho_toggle_block_non_friend_dms = 34
    cho_match_join_success = 36
    cho_match_join_fail = 37
    osu_match_change_slot = 38
    osu_match_ready = 39
    osu_match_lock = 40
    osu_match_change_settings = 41
    cho_fellow_spectator_joined = 42
    cho_fellow_spectator_left = 43
    osu_match_start = 44
    cho_all_players_loaded = 45
    cho_match_start = 46
    osu_match_score_update = 47
    cho_match_score_update = 48
    osu_match_complete = 49
    cho_match_transfer_host = 50
    osu_match_change_mods = 51
    osu_match_load_complete = 52
    cho_match_all_players_loaded = 53
    osu_match_no_beatmap = 54
    osu_match_not_ready = 55
    osu_match_failed = 56
    cho_match_player_failed = 57
    cho_match_complete = 58
    osu_match_has_beatmap = 59
    osu_match_skip_request = 60
    cho_match_skip = 61
    cho_unauthorized = 62  
    osu_channel_join = 63
    cho_channel_join_success = 64
    cho_channel_info = 65
    cho_channel_kick = 66
    cho_channel_auto_join = 67
    osu_beatmap_info_request = 68
    cho_beatmap_info_reply = 69
    osu_match_transfer_host = 70
    cho_privileges = 71
    cho_friends_list = 72
    osu_friend_add = 73
    osu_friend_remove = 74
    cho_protocol_version = 75
    cho_main_menu_icon = 76
    osu_match_change_team = 77
    osu_channel_part = 78
    osu_receive_updates = 79
    cho_monitor = 80  
    cho_match_player_skipped = 81
    osu_set_away_message = 82
    cho_user_presence = 83
    osu_irc_only = 84
    osu_user_stats_request = 85
    cho_restart = 86
    osu_match_invite = 87
    cho_match_invite = 88
    cho_channel_info_end = 89
    osu_match_change_password = 90
    cho_match_change_password = 91
    cho_silence_end = 92
    osu_tournament_match_info_request = 93
    cho_user_silenced = 94
    cho_user_presence_single = 95
    cho_user_presence_bundle = 96
    osu_user_presence_request = 97
    osu_user_presence_request_all = 98
    osu_toggle_block_non_friend_dms = 99
    cho_user_dm_blocked = 100
    cho_target_is_silenced = 101
    cho_version_update_forced = 102
    cho_switch_server = 103
    cho_account_restricted = 104
    cho_rtx = 105 
    cho_match_abort = 106
    cho_switch_tournament_server = 107
    osu_tournament_join_match_channel = 108
    osu_tournament_leave_match_channel = 109
}