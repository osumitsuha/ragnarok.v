module objects

pub struct Match {
	penis	string
}