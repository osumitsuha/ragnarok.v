module managers

pub struct Channel {
	penis	string
}