module constants

const (
	banned 			= 1 << 0

	user 			= 1 << 1
	verified 		= 1 << 2

	supporter 		= 1 << 3

	bat 			= 1 << 4
	moderator 		= 1 << 5
	admin			= 1 << 6
	dev				= 1 << 7

	pending 		= 1 << 8
)