module main
  
const (
    sql_pass  = "password"
    sql_username = "root"
    sql_host = "127.0.0.1"
    sql_table = "ragnarok"

    avatar_domain = "http://127.0.0.1:1001"
    domain = "http://127.0.0.1:1002"
)
