module objects

pub struct Channel {
	penis	string
}