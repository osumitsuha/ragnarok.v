module managers

pub struct Match {
	penis	string
}